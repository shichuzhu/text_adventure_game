{"location":"Cross","inventory":["233-A+","handout","225-A+","I-card","241-A+","I-clicker"],"quests":{"Master-Computer-Science":{"desc":"Take all the three core courses (CS225, CS233, CS241) and then celebrate at home."}},"id":"p0","tick":{"p0":51},"the-map":{"Home":{"desc":"Home, sweet home. No more time for bed because it's a new semester! Before heading out, remember to 'look' around in the room for useful things to bring with you. Use 'quest' to check your goal.","title":"at home","dir":{"north":"Cross"},"contents":[],"events":{"GamePoint":{"hint-text":"'Celebrate' once you completed the three courses.","post-text":"You have finished this game. Congrats! You now master the essence of computer science!","require":["233-A+","225-A+","241-A+"],"match-words":["celebrate"],"questDone":"Master-Computer-Science","action":["[:_configuration] #(assoc % :finished true)"]}}},"Cross":{"desc":"You need to make the hardest decision on which course to take. Choose which building to go. There will be a course available in each of them. Some Easter eggs are on the ground.","title":"at the life's crossroad","dir":{"north":"ECE","south":"Home","west":"DCL","east":"Siebel"},"contents":[]},"Rm1320":{"desc":"You meet Geoffrey here. Get ready for some architecture.","title":"in DCL Rm1320","dir":{"south":"DCL"},"contents":[],"events":{}},"ECE":{"desc":"Good morning\/afternoon! This is cs225. Here is the ECE building. Don't forget to grab a handout.","title":"in the ECE auditorium","dir":{"south":"Cross"},"contents":[],"events":{}},"_quests":{"Master-Computer-Science":{"desc":"Take all the three core courses (CS225, CS233, CS241) and then celebrate at home."},"The-Egg-Hunter":{"desc":"Return the raw-egg to the right hand."},"Data-Structures":{"desc":"cs225 Dear Wade & Mattox!"},"System-Programming":{"desc":"cs241 Threads, pthreads, pppppppp-threads!"},"Architecture":{"desc":"cs233 Spim dat bot!"}},"Rm1304":{"desc":"Welcome to cs241. The creator of the game is lazy -- just sit down and 'learn' the course.","title":"in Siebel Rm1304","dir":{"north":"Siebel"},"contents":[],"events":{}},"_configuration":{"StartingLocation":"Home","StartingQuests":["Master-Computer-Science"],"StartingInventory":[]},"_itemAttr":{"raw-egg":{"desc":"Some poor guy might be desperately looking for his\/her Eastern egg. Oh, Ethan is his name.","questNew":"The-Egg-Hunter"},"I-card":{"desc":"Where there's a card, there's a swiper."},"handout":{"desc":"Quiz today: type any name of the data-structure we learnt this semester to finish this course. Easy, huh?"}},"DCL":{"desc":"Welcome to the Digital Computer Laboratory. Weird as it is, most of the doors are locked inside the building. Some other rooms have card swiper at the door.","title":"in the DCL building","dir":{"east":"Cross","north":"Rm1320"},"contents":[],"events":{}},"Siebel":{"desc":"You've entered the Siebel building. There are a lot people as well as a lot of rooms here. Try to 'talk' to someone asking which is the right room for cs241 here.","title":"in the Siebel Center","dir":{"west":"Cross","south":"Rm1304"},"contents":[],"events":{}}},"seen":["Siebel","Rm1320","Rm1304","Cross","DCL","ECE","Home"]}
